2�d d        d   
 ��  Cand3  ���R  ����                       ��  Cpin  ���  ���0 0                  �  ���  ���0 0                  �  ����  ����1 1                   �Q  ���C  ���0 0                  �  ����S  ����                       �  ����  ����0 0                  �  ����  ����0 0                  �  ����  ����1 1                   �R  ����D  ����0 0                  ��  Cand2  {���S  W���                       �  o���  o���1 1                  �  c���  c���1 1                   �R  i���D  i���1 1                  ��  Cor3�  �����  ����                       ��  �����  ����0 0                  ��  �����  ����0 0                  ��  �����  ����1 1                   ��  �����  ����1 1                  ��  Cswitch   ����)   e���3   ~���L   l��� A    �)   ����)   ����1 0                  �   ����   ����0                     �#   e���#   s���1 0 A    e���        �Z   ����f   f���p   ����   m��� B    �f   ����f   ����1 Z                  �Z   ����Z   ����0                     �`   f���`   t���0 0 B\   f���        ��   �����   f����   ����   m��� C    ��   �����   ����1                    ��   �����   ����0                     ��   f����   t���1 0 C�   f���        ��   �����   e����   ~���
  l��� D    ��   �����   ����1                    ��   �����   ����0                     ��   e����   s���1 0 D�   e���        �� 	 Cinverter   #���[   ����                       �   ���+   ���1 1                   �[   ���M   ���0 0                  )�s   g����   C���                       �s   U����   U���0 0                   ��   U����   U���1 1                  	 ��  Cnet1 	 ��  Csegment#   e���#   e���2�#   e���#   (���2�#   (���   (���2�   ���   (���2�   ���   ���2�   ���   k���2�   k���  k���2�  o���  k���2�  o���  o��� +    0�0  2�`   f���`   ���2�`   f���`   f���2�c   ���  ���2�  ���  ���2�  ���  ���2�`   ���c   ���2�c   ���c   ����2�  ����c   ����2�  ����  ����2�c   ����c   U���2�c   U���s   U���2�s   U���s   U���  
 .    0�1  2��   e����   ����2��   e����   e���2��   ����  ����2�  ����  ����2�  ����  ����   ( 0�0  2�  ���  ���2�[   ���  ���2�[   ���[   ���2�  ���  ���2�[   ���[   ����2�  ����[   ����2�  ����  ����  	  , 0�0  2��  �����  ���2�Q  ����  ���2�Q  ���Q  ���2��  �����  ����    0�0  2�R  �����  ����2�R  ����R  ����2��  �����  ����    0�1  2��  �����  i���2�R  i����  i���2�R  i���R  i���2��  �����  ����    0�1  2��   f����   ����2��   f����   f���2��   ����  ����2�  ����  ����2�  ����  ����   $ 0�1  2�  c���  U���2��   U���  U���2��   U����   U���2�  c���  c���   /   zacharytschirhart