2�d d         d    �� 
 CDflipflop�  i����  ���                       ��  Cpin�  +����  +���1 1                  ��  C����  C���1 1                  ��  i����  [���1 1                  ��  ����  ���1 1                   ��  C����  C���0 0                  ��  +����  +���1 1                  ��  �����  c���                       ��  �����  ����1 1                  ��  �����  ����0 0                  ��  �����  ����1 1                  ��  c����  q���1 1                   ��  �����  ����0 0                  ��  �����  ����1 1                  ��  $����  ����                       ��  �����  ����1 1                  ��  �����  ����0 0                  ��  $����  ���1 1                  ��  �����  ����1 1                   ��  �����  ����0 0                  ��  �����  ����1 1                  ��  Cnand2�   V���.  2���                       ��   J����   J���0 0                  ��   >����   >���1 1                   �-  D���  D���1 1                  ��   �����   ����                       ��   �����   ����1 1                  ��   �����   ����0 0                   ��   �����   ����1 1                  ��   �����   ����                       ��   �����   ����0 0                  ��   �����   ����0 0                   ��   �����   ����1 1                  ��   ����1  ����                       ��   �����   ����1 1                  ��   �����   ����1 1                   �0  ����"  ����0 0                  ��   -����   	���                       ��   !����   !���0 0                  ��   ����   ���1 1                   ��   ����   ���1 1                  ��    ����   ����                       ��   �����   ����0 0                  ��   �����   ����1 1                   ��   �����   ����1 1                  ��   ���6  ����                       ��   ����   ���1 1                  ��   �����   ����1 1                   �5  ���'  ���0 0                  �� 	 CinverterL   �����   ����                       �L   ����Z   ����0 0                   ��   ����|   ����1 1                  5�N   '����   ���                       �N   ���\   ���0 0                   ��   ���~   ���1 1                  5�L   �����   ����                       �L   ����Z   ����0 0                   ��   ����|   ����1 1                  ��  Cprobe:  o���N  O���G  ����a  o���  C     �D  O���D  ]���0 0 C@  O���          ?�>  ����R  ����K  ����d  ����  B     �H  ����H  ����0 0 BD  ����          ?�@  +���T  ���M  =���f  +���  A     �J  ���J  ���0 0 AG  ���          5�P   J����   &���                       �P   8���^   8���0 0                   ��   8����   8���1 1                  ��  Cswitch6  ����B  `���L  y���  g��� Clock    �6  `���6  n���1 0                  �B  `���B  n���0                     �<  ����<  ����1 0 ClockL  y���        I��  �����  ^����  w���<  e��� 	Clear All    ��  ^����  l���1                    ��  ^����  l���0                     ��  �����  ����1 0 	Clear All�  w���        I�W  f����  Z���                       �W  f���e  f���1 0                  �W  Z���e  Z���0                     ��  `���y  `���1 0                  I�^  �����  ����                       �^  ����l  ����1                    �^  ����l  ����0                     ��  �����  ����1 0                  I�^  0����  $���                       �^  0���l  0���1                    �^  $���l  $���0                     ��  *����  *���1 0                   ��  Cnet1  ��  Csegment�  C����  D���`�-  D����  D���`�-  D���-  D���`��  C����  C���    ^�0  `�D  O���D  C���`��  C���D  C���`��  C����  C���`�D  O���D  O���`��  C����  C���`��  C����  }���`��   }����  }���`��   }����   J���`��   J����   J���`��   J����   J���`�   }����   }���`�L   ����L   ����`�   ����   %���`�   %����   %���`��   !����   %���`��   !����   !���`�   %���   ����`�L   ����   ����`�L   ����L   ����`�   ����L   ����`�   ����   }���`�   ����   ���� A  7 * =   ^�0  `�H  ����H  ����`�  ����H  ����`��  �����  ����`�H  ����H  ����`��  ����  ����`�  ����  ����`�8   ����  ����`�8   ����8   8���`�P   8���8   8���`�P   8���P   8���`�8   ����8   ����`�8   �����   ����`��   �����   ����`��   �����   ���� C G "   ^�0  `�J  ���J  ����`�  ����J  ����`��  �����  ����`�J  ���J  ���`��  ����  ����`�  ����  ]���`�B   ]���  ]���`�   ]���   ����`�\   ����   ����`��   �����   ����`��   ����\   ����`�\   ����\   ����`��   ����\   ����`��   �����   ����`�   ]���B   ]���`�B   ]���B   ���`�N   ���B   ���`�N   ���N   ���`�B   ���B   ����`��   ����B   ����`��   �����   ���� E  # : .   ^�1  `��   >����   8���`��   8����   8���`��   8����   8���`��   >����   >���   H ^�1  `��   �����   ����`��   �����   ����`��   �����   ����`��   �����   ����   8 ^�1  `��   �����   ����`��   �����   ����`��   �����   ����`��   �����   ���� &    ^�1  `��   �����   ����`��   �����   ����`��   �����   ����`��   �����   ���� '  $ ^�0  `��  �����  ����`�0  �����  ����`�0  ����0  ����`��  �����  ����   ( ^�1  `��   �����   ����`��   �����   ����`��   �����   ����`��   �����   ���� /  > ^�1  `��   ����   ���`��   ����   ���`��   ����   ��� +  ; ^�1  `��   ����   ���`��   ����   ���`��   ����   ���`��   ����   ��� 2  , ^�1  `��   �����   ����`��   �����   ����`��   �����   ����`��   �����   ���� 3  0 ^�0  `��  �����  ���`�5  ����  ���`�5  ���5  ���`��  �����  ����   4 ^�1 
 `��  ����  ���`��  ����  ���`��  �����  ����`��  c����  c���`��  c����  c���`��  �����  ����`��  �����  ����`��  �����  ����`��  c����  ����`��  c����  ���     Q ^�1 
 `�<  �����  ����`��  �����  ����`�<  ����<  ����`�<  ����<  ����`�<  ����<  ����`��  ����<  ����`��  �����  ����`�<  ����<  +���`��  +���<  +���`��  +����  +���     M ^�1  `��  `����  i���`��  i����  i���`��  i����  i���`��  `����  `���   U ^�1  `��  �����  ����`��  �����  ����`��  �����  ����`��  �����  ����   Y ^�1  `��  *����  $���`��  $����  $���`��  $����  $���`��  *����  *���   ]   zacharytschirhart