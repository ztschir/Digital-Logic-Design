2�d d        d    ��  Cnand3  S���N  /���                       ��  Cpin  M���  M���0 0                  �  A���  A���1 1 D�   O���        �  5���  5���0 0 E'�   C���         �M  A���?  A���1 1 (A'DE')'M  O���        �  ����N  ����                       �  ����  ����0 0 B�   ����        �  ����  ����1 1 D�   ����        �  ����  ����0 0 E'�   ����         �M  ����?  ����1 1 (BDE')'M  ����        ��   b���J  >���                       ��   \���  \���0 0                  ��   P���  P���0 0 D'�   ^���        ��   D���  D���1 1 E�   R���         �I  P���;  P���1 1 (A'D'E)'I  ^���        �  ����M  ~���                       �  ����  ����1 1 B'�   ����        �  ����  ����1 1 D�   ����        �  ����  ����1 1 E�   ����         �L  ����>  ����0 0 (B'DE)'L  ����        ��  Cnand2�   ����E  a���                       ��   y���  y���0 0 B�   ����        ��   m���  m���1 1 E�   {���         �D  s���6  s���1 1 (BE)'D  ����        ��  Cnand48  �����  ����E  ����]  ���� Z     �8  ����F  ����0 0 (AC)'  ����        �8  ����F  ����1 1 (BE)'  ����        �8  ����F  ����1 1 (BCD)'  ����        �8  ����F  ����0 0 (AE)'  ����         ��  ����t  ����1 1 Z�  ����        ��  Cswitch   ����'   w���1   ����J   ~��� A    �'   ����'   ����1 Z                  �   ����   ����0 Z                   �!   w���!   ����1 0 A1   ����        #�F   ����R   y���\   ����u   ���� B    �R   ����R   ����1                    �F   ����F   ����0                     �L   y���L   ����0 0 B\   ����        #�n   ����z   y����   �����   ���� C    �z   ����z   ����1                    �n   ����n   ����0                     �t   y���t   ����1 0 C�   ����        #��   �����   x����   �����   ��� D    ��   �����   ����1                    ��   �����   ����0                     ��   x����   ����1 0 D�   ����        #��   �����   w����   �����   ~��� E    ��   �����   ����1                    ��   �����   ����0                     ��   w����   ����1 0 E�   ����        �� 	 Cinverter   t���>   6���                      �,   t���,   f���1 1                   �,   6���,   D���0 0                  8�:   0���^   ����                      �L   0���L   "���0 0                   �L   ����L    ���1 1 B'G   ����        8�b   0����   ����                      �t   0���t   "���1 1                   �t   ����t    ���0 0 C'o   ����        8��   0����   ����                      ��   0����   "���1 1                   ��   �����    ���0 0 D'�   ����        8��   0����   ����                      ��   0����   "���1 1                   ��   �����    ���0 0 E'�   ����        �>  ]����  9���                       �>  Q���L  Q���1 1                  �>  E���L  E���1 1 D.  I���         ��  K���z  K���0 0 (AD)'�  Y���        �=  ����  ����                       �=  	���K  	���0 0 B5  ���        �=  ����K  ����1 1 D4  ���        �=  ����K  ����1 1 E5  ����         ��  ����y  ����1 1 (BDE)'�  ���        �(  <���s  ���5  N���R  <��� W     �(  6���6  6���0 0 (AD)'  D���        �(  *���6  *���0 0 C'  8���        �(  ���6  ���1 1 (BDE)'  ,���         �r  *���d  *���1 1 Wr  8���        ��  Cnand5-  ����x  b���:  ����R  ���� X     �-  ����;  ����1 1 (A'DE')'  ����        �-  ����;  ����1 1 (BC)'  ����        �-  u���;  u���0 0 (B'DE)'  ����        �-  i���;  i���0 0 (AE)'  w���        �-  ]���;  ]���0 0 (AC)'  k���         �w  t���i  t���1 1 Xw  ����        �%  ����p  w���                       �%  ����3  ����0 0 B  ����        �%  ����3  ����1 1 C  ����         �o  ����a  ����1 1 (BC)'o  ����        ��  0����  ���                       ��  $����  $���1 1 A�  2���        ��  ����  ���1 1 E�  &���         ��  ����  ���0 0 (AE)'�  ,���        ��  �����  ����                       ��  �����  ����1 1 A�   ���        ��  �����  ����1 1 C�  ����         ��  �����  ����0 0 (AC)'�  ����        V�D  N����  *���Q  `���j  N��� Y     �D  U���R  U���0 0                  �D  I���R  I���0 0 (AC)'*  W���        �D  =���R  =���0 0 (AD)'*  K���        �D  1���R  1���0 0 (CE)')  ?���        �D  %���R  %���1 1 (BDE')'!  3���         ��  <����  <���1 1 Y�  J���        ��  Cand2�  y���C  U���                       ��  m���  m���1 1 (A'D'E)'�  {���        ��  a���  a���0 0 (B'DE)'�  o���         �B  g���4  g���0 0                  �  ����L  ����                       �  ����  ����1 1 C�   ����        �  ����  ����1 1 E�   ����         �K  ����=  ����0 0 (CE)'K  ����        ��   ����J  ����                       ��   ����  ����0 0 B�   ����        ��   ����  ����1 1 C�   ����        ��   ����  ����1 1 D�   ����         �I  ����;  ����1 1 (BCD)'I  ����        ��  Cprobe�  S����  3���                        ��  3����  A���1 1                    ��  U����  5���                        ��  5����  C���1 1                    ��  U����  5���                        ��  5����  C���1 1                    ��  U����  5���                        ��  5����  C���1 1                    # ��  Cnet0      ' ��0  ��  CsegmentL   0���L   0�����L   0���L   y�����L   y���L   y��� = 	  M _ {  + ��1  ���   0����   0������   0����   x������   x����   x������   x����   x��� C J  
  N }  3 ��0    S  A ��Z  ��>  I���>  J���    ��Z       ��Z       ��Z       ��Z       ��1  ��,   t���,   t�����!   t���,   t�����!   w���!   w�����!   w���!   �������   ����  ������  w���  ������>  w���  w�����>  Q���>  Q�����!   �����   �������   �����   �����   ����   �����>  Q���>  w�����   ���   $������  $���   $������  $����  $�����   ����  ������  �����  ������  �����  ������!   t���!   ���� : I c g  ' ��0 
 ��@   6���V   6�����V   ����V   6�����,   6���,   6�����  M���  ������  M���  M�����,   6���@   6�����@   6���@   \������   \���@   \������   \����   \�����V   ����  ����    ; ��0       G ��1      > ��0      D ��Z  ��2  9���2  :���    ��1  ��t   0���t   0�����t   y���t   0�����t   y���t   y��� @ ` h w |  / ��Z       ��0    R m  K ��1    T  P ��1    X   ��1    Y  a ��0    [ !  e ��0    \ l   i ��0    Z t   ��0  ��B  g���B  g�����D  U���D  U�����D  g���B  g�����D  U���D  g��� k  u ��1    s   ��0    n  y ��1       ��1  ���  3����  *�����r  *����  *�����r  *���r  *������  3����  3��� �  U ��1  ���  5����  t�����w  t����  t�����w  t���w  t������  5����  5��� �  ] ��1  ���  5����  <������  <����  <������  <����  <������  5����  5��� �  p ��1  ���  5����  �������  �����  �������  �����  �������  5����  5��� �  " ��1    o   ��1  ���   0����   0������   0����   w������   w����   w������   w����   w��� F    O d x  7 ��1  ��8  ����8  ������8  ����8  ����    ~   zacharytschirhart