2�d d         d     ��  Cnor3  {���S  W���                       ��  Cpin  u���  u���1 1                  �  i���  i���0 0 B   w���        �  ]���  ]���1 1 C�   k���         �R  i���D  i���0 0                  �	  ���T  ����                       �	  ���  ���1 1 B'�   ���        �	  ����  ����1 1 C   ���        �	  ����  ����1 1 E  ����         �S  ����E  ����0 0                  ��  Cnor2	  A���T  ���                       �	  5���  5���1 1 C   C���        �	  )���  )���1 1 D   7���         �S  /���E  /���0 0                  ��  A���  ���                       ��  ;����  ;���0 0                  ��  /����  /���0 0                  ��  #����  #���0 0                   �  /����  /���1 1 W  =���        ��  Cswitch"   ����.   ����%   ����>   ���� A    �.   ����.   ����1 0                  �"   ����"   ����0 Z                   �(   ����(   ����1 0 A%   ����        �G   ����S   ����I   ����b   ���� B    �S   ����S   ����1 Z                  �G   ����G   ����0                     �M   ����M   ����0 0 BI   ����        �r   ����~   ����t   �����   ���� C    �~   ����~   ����1                    �r   ����r   ����0                     �x   ����x   ����1 0 Ct   ����        ��   �����   �����   �����   ���� D    ��   �����   ����1                    ��   �����   ����0                     ��   �����   ����1 0 D�   ����        ��   �����   �����   �����   ���� E    ��   �����   ����1                    ��   �����   ����0                     ��   �����   ����1 0 E�   ����        �� 	 Cinverter   ����<   ����                      �*   ����*   ����1 1                   �*   ����*   ����0 0 A'&   ����        ,�=   p���a   2���                      �O   p���O   b���0 0                   �O   2���O   @���1 1 B'J   2���        ,�e   q����   3���                      �w   q���w   c���1 1                   �w   3���w   A���0 0 C'r   3���        ,��   q����   3���                      ��   q����   c���1 1                   ��   3����   A���0 0 D'�   3���        ,��   p����   2���                      ��   p����   b���1 1                   ��   2����   @���0 0 E'�   2���        �
  ����U  ����                       �
  ����  ����1 1                  �
  ����  ����0 0 B  ����        �
  ����  ����1 1 D  ����         �T  ����F  ����0 0                  �  ����S  w���                       �  ����  ����1 1 B'�   ����        �  ����  ����1 1 C�   ����        �  }���  }���0 0 E'�   ����         �R  ����D  ����0 0                  �  l���P  H���                       �  f���  f���0 0                  �  Z���  Z���1 1 C�   h���        �  N���  N���1 1 E�   \���         �O  Z���A  Z���0 0                  �  A���R  ���                       �  ;���  ;���1 1 B'�   I���        �  /���  /���1 1 C�   =���        �  #���  #���1 1 D�   1���         �Q  /���C  /���0 0                  ��  Cnor4�  ����
  c���                       ��  �����  ����0 0                  ��  {����  {���0 0                  ��  o����  o���0 0                  ��  c����  c���0 0                   �	  u����  u���1 1 X	  ����        �  ���S  ����                       �  ���  ���1 1                  �  ���  ���0 0 B   ���        �  ����  ����1 1 E   ���         �R  ���D  ���0 0                  �	  ����T  ����                       �	  ����  ����0 0                  �	  ����  ����1 1 C   ����        �	  ����  ����1 1 D   ����         �S  ����E  ����0 0                  �  |���R  X���                       �  v���  v���1 1 B'�   ����        �  j���  j���1 1 D�   x���        �  ^���  ^���1 1 E�   l���         �Q  j���C  j���0 0                  P�	  ����T  ����                       �	  ����  ����1 1 B'�   ����        �	  ����  ����1 1 C   ����        �	  ����  ����0 0 D'�   ����        �	  ����  ����0 0 E'�   ����         �S  ����E  ����0 0                  P��  �����  ����                       ��  �����  ����0 0                  ��  �����  ����0 0                  ��  �����  ����0 0                  ��  �����  ����0 0                   ��  �����  ����1 1 Y�  ����        �  E���R  !���                       �  9���  9���1 1                  �  -���  -���0 0 B�   ;���         �Q  3���C  3���0 0                  �  ���R  ����                       �  ���  ���1 1 C�   ���        �   ���   ���1 1 E�   ���         �Q  ���C  ���0 0                  �  ����S  ����                       �  ����  ����1 1 B'�   ����        �  ����  ����1 1 D�   ����        �  ����  ����1 1 E   ����         �R  ����D  ����0 0                  ��  ����  ����                       ��  ����  ���0 0                  ��  ����  ���0 0                  ��  �����  ����0 0                   ��  ����  ���1 1 Z�  ���        ��  Cprobe/  ����C  n���                        �9  n���9  |���1 1                    ��H  ����\  o���                        �R  o���R  }���1 1                    ��b  ����v  o���                        �l  o���l  }���1 1                    ��|  �����  o���                        ��  o����  }���1 1                     ��  Cnet1  ��  Csegment*   ���*   ������(   ����*   ������(   ����(   ������*   ����*   ������*   ����*   �����*   ����   ������   u����   ������   u���  u�����  u���  u������   �����   �����
  ����
  �������   ����   ������  ���  �����
  �����   ������  ����   ������   ����   9�����  9����   9�����  9���  9��� .  = X s   ��0  ��O   p���O   ������M   ����O   ������M   ����M   ������O   p���O   p��� 1  > Y t   ��1  ��w   q���w   ������x   ����w   ������x   ����x   ������w   q���w   q���
 4   
 C H M ^ h w  # ��1  ���   �����   q������   �����   �������   q����   q��� 7  ? N _ c |  ' ��1  ���   p����   �������   �����   �������   �����   �������   p����   p��� :  I Z d x }  + ��1    	 B L g b {  2 ��0  ���  i���R  i�����R  i���R  i������  ;����  ;������  ;����  i���    ��0  ��S  /���S  /������  /����  /������  /���S  /���    ��0  ���  ����S  ������S  ����S  �������  #����  #������  #����  ����    ��0  ��*   f���*   ������*   ����*   ������  f���  f�����*   ����*   f�����	  ����	  ������  f���*   f�����	  ����*   ���� G ]  / ��0    D j  ; ��0  ��T  ����T  �������  �����  �������  ����T  �������  �����  ���� R  @ ��0  ��R  ����R  ������T  ����R  ������T  {����  {������  {����  {�����T  ����T  {��� S  E ��0  ��O  Z���O  Z������  o����  o�����U  o����  o�����U  Z���O  Z�����U  o���U  Z��� T  J ��0  ��Q  /���Q  /������  c����  c������  /���Q  /������  c����  /��� U  O ��0    i  8 ��0  ���  �����  �����R  ����  �����R  ���R  ������  �����  ���� m  [ ��0  ��S  �����  �������  �����  ������S  ����S  �������  �����  �������  �����  �������  �����  ���� n  ` ��0  ��S  ����~  ������~  ����~  ������S  ����S  ������~  �����  �������  �����  �������  �����  ���� o  k ��0  ���  �����  j�����Q  j����  j�����Q  j���Q  j������  �����  ���� p  e ��0  ���  ����  3�����Q  3����  3�����Q  3���Q  3������  ����  ��� �  u ��0  ��Q  ����  �����Q  ���Q  ������  ����  ��� �  y ��0  ���  �����  ������R  �����  ������R  ����R  �������  �����  ���� �  ~ ��1  ��9  n���9  /�����  /���9  /�����  /���  /�����9  n���9  n��� �   ��1  ��R  o���R  u�����	  u���R  u�����	  u���	  u�����R  o���R  o��� �  V ��1  ��l  o���l  �������  ����l  �������  �����  ������l  o���l  o��� �  q ��1  ���  o����  ������  ����  ������  ����  ������  o����  o��� �  �   zst75