5�d d         �	   �� 
 CDflipflope  9����  ����                       ��  Cpine  ����s  ����0 0                  �e  ���s  ���0 0                  ��  9����  +���1 1                  ��  �����  ����0 0                   ��  ����  ���0 0 Q1�  !���        ��  �����  ����1 1 Q1'�  	���        �f  �����  N���                       �f  t���t  t���0 0                  �f  ����t  ����1 1                  ��  �����  ����1 1                  ��  N����  \���0 0                   ��  �����  ����0 0 Q2�  ����        ��  t����  t���1 1 Q2'�  ����        �f  &����  ����                       �f  ����t  ����0 0                  �f   ���t   ���1 1                  ��  &����  ���Z Z                  ��  �����  ����0 0                   ��   ����   ���0 0 Q3�  ���        ��  �����  ����1 1 Q3'�  ����        ��  Cnand2�   ���G  ����                       ��   ���
  ���1 1                  ��   ����
  ����0 0 X�   ���         �F  ����8  ����1 1                  �m   �����   q���                       �m   ����{   ����0 0 Q1]   ����        �m   }���{   }���0 0 Q3]   ����         ��   �����   ����1 1                  ��   ;����   ���                       ��   /����   /���0 0 Q3�   =���        ��   #����   #���1 1 X'�   1���         ��   )����   )���1 1                  ��   ����   ����                       ��   �����   ����1 1 Q2'�   	���        ��   �����   ����0 0 Q3�   ����         ��   �����   ����1 1                  ��  Cnand3  "���X  ����                       �  ���  ���1 1                  �  ���  ���1 1                  �  ���  ���1 1                   �W  ���I  ���0 0                  )��   o���A  K���                       ��   i���  i���0 0 Q2�   w���        ��   ]���  ]���1 1 X'�   k���        ��   Q���  Q���1 1 Q3'�   _���         �@  ]���2  ]���1 1                  ��  Cnor3  ����d  m���                       �  ����,  ����1 1                  �  ���-  ���0 0                  �  s���,  s���0 0 X  ����         �c  ���U  ���0 0 Zc  ����        ��  Cprobex  �����  ����  �����  o���  Z     ��  �����  ����0 0 Z  ����          �� 	 Cinverter^  �����  ����                      �p  ����p  ����0 0                   �p  ����p  ����1 1 X'l  ����        :�  ����1  ����  ����B  p���  Q1     �'  ����'  ����0 0 Q1  ����          :�9  ����M  ����;  ����^  q���  Q2     �C  ����C  ����0 0 Q2;  ����          :�T  ����h  ����W  ����z  s���  Q3     �^  ����^  ����0 0 Q3W  ����          ��  CplusV�  �����  ����                          ��  �����  ����1 1                  G��  �����  ����                          ��  �����  ����1 1                  G��  �����  ����                          ��  �����  ����1 1                  ��  Cswitch�  �����  ^����  �����  ���� rst    ��  ^����  l���1 0                  ��  ^����  l���0 1                   ��  �����  ����0 0 rst�  ����        N�0  S���<  #���F  <���^  *��� X    �0  #���0  1���1 1                  �<  #���<  1���0 ��                  �6  S���6  E���0 0 X3  a���        N�  C���?  7���  U���=  C��� clk     �  C���  C���1 1                  �  7���  7���0                     �?  =���1  =���0 0 clk?  K���         ��  Cnet1  ��  Csegment  ���  )���]��   )���  )���]��   )����   )���]�  ���  ��� +  $ [�1  ]��   �����   ����]��   ����   ����]��   �����   ����]��   ���  ���]�  ���  ���]�  ���  ���]�  ���  ��� ,  ( [�1 	 ]��   �����   ����]��   �����   ����]��   �����   ����]��   ����  ����]�  ���  ����]�  ���  ���]��   �����   ���]��   ����   ���]��   ����   ��� -     [�1  ]�@  ]���F  ]���]�F  ����F  ]���]�@  ]���@  ]���]�F  ����f  ����]�f  ����f  ����]�f  ����f  ����   3 [�1  ]�  ����  ����]��  ����  ����]��  �����  ����]�  ����  ���� 6  	 [�1  ]�F  ����F   ���]�f   ���F   ���]�f   ���f   ���]�F  ����F  ����    [�0  ]�e  ���e  ���]�W  ���e  ���]�W  ���W  ���]�e  ���e  ���   . [�0  ]��  ���c  ���]�c  ���c  ���]��  �����  ����]��  ����  ���� <  9 [�0  ]��  N����  ����]��  �����  ����]��  �����  ����]��  N����  N���]��  �����  N���]��  N����  N���]��  �����  ����]��  �����  ����]��  �����  ����]��  ~����  ����]��  �����  ����]��  �����  ����]��  �����  ����     R [�0  ]�p  ����p  ����]�p  ����p  }���]�3  k���3  }���]�3  }���p  }���]�3  `���3  k���]�6  k���3  k���]�6  S���6  k���]�6  S���6  S���  8 ?  V [�1  ]��  9����  ����]��  9����  9���]��  �����  ����]��  �����  ����]��  �����  ����   I [�1  ]��  �����  ����]��  �����  ����]��  �����  ����]��  �����  ����]��  �����  ����]��  �����  ����]��  �����  ����]��  �����  ����   K [�1    # 1  @ [�Z  �     [�1  ]��  |����  !���]��  !����  !���]��  �����  |���]��  |����  |���]��  �����  |���]��  �����  ����   M [�Z       [�0  ]�e  ����e  ����]�e  ����_  ����]�_  t���_  ����]�_  t���f  t���]�_  ����_  t���]�_  ����f  ����]�_  ?���_  ����]�f  ����f  ����]�f  t���f  t���]�_  <���_  ?���]�_  ?���?  ?���]�?  =���?  ?���]�?  =���?  =���     Z [�Z       [�1    2   [�0  ]�C  ����C  ����]�C  ����A  ����]�A  	���A  ����]�A  	���  	���]�  ����  	���]��  ����  ����]��  �����  ���� D 0   [�Z  ]�'  ����'  ����]�'  ����'  ���]��  ���'  ���]��  ����  ��� B    [�0 
 ]�  ���  ���]�  ���  ~���]��  ~���  ~���]��  ~����   ���]��   ����   ���]�_   ����   ���]�_   ���_  ����]�^  ����_  ����]�^  ����^  ����]��   ����   ��� 7 F  " '   [�1    &     zst75