5�d d       �	   ��  Cclock  E���7  3���                2         ��  Cpin7  <���)  <���0 1                  �� 
 CDflipflope  9����  ����                       �e  ����s  ����0 0                  �e  ���s  ���1 1                  ��  9����  +���1 1                  ��  �����  ����1 1                   ��  ����  ���1 1 Da�  !���        ��  �����  ����0 0 Da'�  	���        �f  �����  N���                       �f  t���t  t���0 0                  �f  ����t  ����1 1                  ��  �����  ����1 1                  ��  N����  \���1 1                   ��  �����  ����1 1 Db�  ����        ��  t����  t���0 0 Db'�  ����        �f  &����  ����                       �f  ����t  ����0 0                  �f   ���t   ���1 1                  ��  &����  ���1 1                  ��  �����  ����1 1                   ��   ����   ���1 1 Dc�  ���        ��  �����  ����0 0 Dc'�  ����        ��  Cnand2�   ���G  ����                       ��   ���
  ���0 0                  ��   ����
  ����0 0 X�   ���         �F  ����8  ����1 1                  �m   �����   q���                       �m   ����{   ����1 1 Da]   ����        �m   }���{   }���1 1 Dc^   ����         ��   �����   ����0 0                  ��   ;����   ���                       ��   /����   /���1 1 Dc�   =���        ��   #����   #���1 1 X'�   1���         ��   )����   )���0 0                  ��   ����   ����                       ��   �����   ����0 0 Db'�   	���        ��   �����   ����1 1 Dc�   ����         ��   �����   ����1 1                  ��  Cnand3  "���X  ����                       �  ���  ���0 0                  �  ���  ���1 1                  �  ���  ���0 0                   �W  ���I  ���1 1                  ,��   o���A  K���                       ��   i���  i���1 1 Db�   w���        ��   ]���  ]���1 1 X'�   k���        ��   Q���  Q���0 0 Dc'�   _���         �@  ]���2  ]���1 1                  ��  Cnor3  ����d  m���                       �  ����,  ����0 0                  �  ���-  ���1 1                  �  s���,  s���0 0 X  ����         �c  ���U  ���0 0 Zc  ����        ��  Cprobex  �����  ����  �����  o���  Z     ��  �����  ����0 0 Z  ����          �� 	 Cinverter^  �����  ����                      �p  ����p  ����0 0                   �p  ����p  ����1 1 X'l  ����        ��  Cswitchd  ����p  ����]  �����  s��� PreA    �p  ����p  ����1 0                  �d  ����d  ����0                     �j  ����j  ����1 1 PreA]  ����        D��  �����  �����  �����  s��� PreB    ��  �����  ����1                    ��  �����  ����0                     ��  �����  ����1 1 PreB�  ����        D��  �����  �����  �����  r��� PreC    ��  �����  ����1                    ��  �����  ����0 ��                  ��  �����  ����1 1 PreC�  ����        =�  ����3  ����,  ����_  ����  Clock     �)  ����)  ����0 0 Clock  ����          =�A  ����U  ����H  ����`  ����  X     �K  ����K  ����0 0 XH  ����          ��  Cchecker�  I���$  ����                       ��   ����   ���0 0                  ��  �����  ���0 0                   ��  I����  ;���1 1                  �$   ���   ���0 0                  101011101001R010101001010000100000100X000010100000 ��  Cnet0  ��  Csegment  ���  )���]��   )���  )���]��   )����   )���]�  ���  ��� .  ' [�1  ]��   �����   ����]��   ����   ����]��   �����   ����]��   ���  ���]�  ���  ���]�  ���  ���]�  ���  ��� /  + [�0 	 ]��   �����   ����]��   �����   ����]��   �����   ����]��   ����  ����]�  ���  ����]�  ���  ���]��   �����   ���]��   ����   ���]��   ����   ��� 0   # [�1  ]�@  ]���F  ]���]�F  ����F  ]���]�@  ]���@  ]���]�F  ����f  ����]�f  ����f  ����]�f  ����f  ����   6 [�0  ]�  ����  ����]��  ����  ����]��  �����  ����]�  ����  ���� 9   [�1  ]�  ���  ���]�  ���  ~���]��  ~���  ~���]��  ~����   ���]��   ����   ���]��   ����   ��� : % * "   [�1  ]�F  ����F   ���]�f   ���F   ���]�f   ���f   ���]�F  ����F  ����    [�0    )   [�1    !   [�1  ]��  �����  ����]��  ����  ���� 3   [�0    5   [�1  ]�e  ���e  ���]�W  ���e  ���]�W  ���W  ���]�e  ���e  ���   1 [�0  ]��  ���c  ���]�c  ���c  ���]��  �����  ����]��  �����  ���]��  �����  ����]��  �����  ����]��   ����  ����]��   ����   ��� ? W  < [�1  ]��  N����  ����]��  �����  ����]��  �����  ����]��  N����  N���]��  �����  N���]��  N����  N���]��  �����  ����]��  �����  ����]��  �����  ����]��  ~����  ����]�  �����  ����]��  I���  I���]�  ����  I���]��  I����  I��� 
    Y [�0  ]�_  t���_  ����]�e  ����_  ����]�e  ����e  ����]�_  t���f  t���]�_  ����_  t���]�f  t���f  t���]�_  ����f  ����]�_  ����_  ����]�f  ����f  ����]�_  ����)  ����]�_  <���_  ����]�)  ����)  ����]�7  <���7  <���]�B  <���_  <���]�7  <���B  <���]�B  3���B  <���]�%  �����  ����]��  �����  ����]�%  H���%  ����]��  3���B  3���]��  H���%  H���]��  H����  3���    R X   [�0  ]�p  ����p  ����]�p  ����p  }���]�K  }���p  }���]�3  }���K  }���]�K  }���K  ����]�K  ����K  ����]�3  `���3  }���]�3  `���V  `���]�V  !���V  `���]�V  !���$  !���]�$   ���$  !���]�$   ���$   ��� B T ;   Z [�1  ]��  9����  ����]�j  �����  ����]�j  ����j  ����]��  9����  9��� 	  H [�1  ]��  �����  ����]��  �����  ����]��  �����  ����]��  �����  ����]��  �����  ����]��  �����  ����   L [�1  ]��  �����  !���]��  �����  ����]��  !����  !���]��  &����  !���]��  &����  &���   P [�1    4 &  C   zst75